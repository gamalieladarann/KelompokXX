module dev(
    input wire signed [19:0] D_out, // Input from var module

    output wire signed [19:0] S_out // Output from dev module
);